// Henry Heathwood
// hheathwood@Hmc.edu
// 9/3/24
// Top level verilog file for lab 1